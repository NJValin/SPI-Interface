/////////////////////////////////////////////////////////////////
// Copyright (c) 2025 Neil Valin. All Rights Reserved.
//
//
/////////////////////////////////////////////////////////////////

`default_nettype none

module spi_top #(
	parameter DATA_WIDTH   = 8,
	parameter BUFFER_DEPTH = 4,
	parameter MASTER = 0       // Determines if the SPI interface will act as a master or a slave
	)
	(
	input  logic                  clk, // Will be gated to form sclk
	input  logic [DATA_WIDTH-1:0] data_in,
	output logic [DATA_WIDTH-1:0] data_out,

	input  logic                   write,
	input  logic                   read,

	// CSR values. The associated registers should be generated by integrating project
	input  logic                  enable,       //SPI enable
	input  logic                  spi_3wire,    // If set, mosi will be used for both read and write transactions
	input  logic                  stop_in_idle, // Stop in IDLE mode
	input  logic                  cpol,         // Clock polarity in IDLE mode
	input  logic                  cpha,         // determines clock phase
	input  logic                  msb_first,    // If set, the msb will be shifted out first, else lsb will be first
	output logic				  rx_v,         // Overflow in receiving flag
	output logic                  tx_buf_full,  // Transmit buffer full
	output logic                  rx_buf_full,  // Receive buffer full


	inout  tri                    cs_b,
	inout  tri                    mosi,
	inout  tri                    miso,
	inout  tri                    sclk
	);

	generate
		if (MASTER==1) begin : MASTER_INTERFACE
			logic                         master_CS_b;
			logic                         master_clock;
		end
		else begin : SLAVE_INTERFACE
			
		end
	endgenerate
	logic                         in_idle;

	assign CS_b = (MASTER==1'b1)?master_CS_b:1'bz; // In slave mode, the value resolved will be the val driven by the master
	
	
endmodule
